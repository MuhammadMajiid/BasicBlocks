module VedicMul_8x8
(
    input wire [7:0] multiplicand,
    input wire [7:0] multiplier,

    output wire [15:0] result
);


    
endmodule